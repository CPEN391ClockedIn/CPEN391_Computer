LIBRARY 	ieee  ;
USE		ieee.std_logic_1164.all ;
use 		IEEE.numeric_std.all;  


----------------------------------------------------------------------------------
-- Top level WHOLE system not just Qsys generated HPS component
----------------------------------------------------------------------------------

entity MyComputer is
	PORT (
		---------------------------------------------
		-- FPGA Pins
		---------------------------------------------
	
		-- Clock pins
		CLOCK_50,CLOCK2_50,CLOCK3_50,CLOCK4_50		: in std_logic; 
		
		-- Seven Segment Displays
		-- These are the names of the 6 seven segment display on the DE1 and those in the PIN Planner,
		--	so stick to these names.
		HEX0,HEX1,HEX2,HEX3,HEX4,HEX5 : out std_logic_vector(6 downto 0) ;
	
		-- Pushbuttons
		KEY			: in std_logic_vector(3 downto 0);
	
		-- LEDs
		LEDR			: out std_logic_vector(9 downto 0);
	
		-- Slider Switches
		SW				: in std_logic_vector(9 downto 0);
		
		-- VGA/Graphics Signals
		VGA_BLANK_N 	:  OUT  STD_LOGIC;
		VGA_SYNC_N		:  OUT STD_LOGIC ;
		
		VGA_CLK 			:  OUT  STD_LOGIC;
		VGA_HS 			:  OUT  STD_LOGIC;
		VGA_VS 			:  OUT  STD_LOGIC;
		
		VGA_B 			:  OUT  STD_LOGIC_VECTOR(7 DOWNTO 0);
		VGA_G 			:  OUT  STD_LOGIC_VECTOR(7 DOWNTO 0);
		VGA_R 			:  OUT  STD_LOGIC_VECTOR(7 DOWNTO 0);
		
	
		-- SDRAM on FPGA Side
		DRAM_ADDR		: out std_logic_vector(12 downto 0);
		DRAM_BA			: out std_logic_vector(1 downto 0);
		DRAM_CAS_N		: out std_logic ;
		DRAM_CKE			: out std_logic ;
		DRAM_CLK			: out std_logic ;
		DRAM_CS_N		: out std_logic ;
		DRAM_DQ			: inout std_logic_vector(15 downto 0);
		DRAM_LDQM		: out std_logic ;
		DRAM_RAS_N		: out std_logic ;
		DRAM_UDQM		: out std_logic ;
		DRAM_WE_N		: out std_logic ;
		
		-- 40-Pin Headers
		GPIO_0			: inout std_logic_vector(35 downto 0);
		GPIO_1			: inout std_logic_vector(35 downto 0);
		

		------------------------------------------------------
		-- HPS Pins
		------------------------------------------------------
		
		-- DDR3 SDRAM
		HPS_DDR3_ADDR		: out std_logic_vector(14 downto 0);
		HPS_DDR3_BA			: out std_logic_vector(2 downto 0);
		HPS_DDR3_CAS_N		: out std_logic ;
		HPS_DDR3_CKE		: out std_logic ;
		HPS_DDR3_CK_N		: out std_logic ;
		HPS_DDR3_CK_P		: out std_logic ;
		HPS_DDR3_CS_N		: out std_logic ;
		HPS_DDR3_DM			: out std_logic_vector(3 downto 0);
		HPS_DDR3_DQ			: inout std_logic_vector(31 downto 0);
		HPS_DDR3_DQS_N		: inout std_logic_vector(3 downto 0);
		HPS_DDR3_DQS_P		: inout std_logic_vector(3 downto 0);
		HPS_DDR3_ODT		: out std_logic ;
		HPS_DDR3_RAS_N		: out std_logic ;
		HPS_DDR3_RESET_N	: out std_logic ;
		HPS_DDR3_RZQ		: in std_logic ;
		HPS_DDR3_WE_N		: out std_logic ;
		
		-- Ethernet
		HPS_ENET_GTX_CLK	: out std_logic ;	
		HPS_ENET_INT_N		: inout std_logic ;
		HPS_ENET_MDC		: out std_logic ;
		HPS_ENET_MDIO		: inout std_logic ;
		HPS_ENET_RX_CLK	: in std_logic;
		HPS_ENET_RX_DATA	: in std_logic_vector(3 downto 0);
		HPS_ENET_RX_DV		: in std_logic;
		HPS_ENET_TX_DATA	: out std_logic_vector(3 downto 0);
		HPS_ENET_TX_EN		: out std_logic ;
	
		-- Flash
		HPS_FLASH_DATA		: inout std_logic_vector(3 downto 0);
		HPS_FLASH_DCLK		: out std_logic ;	
		HPS_FLASH_NCSO		: out std_logic ;	
	
		-- Accelerometer
		HPS_GSENSOR_INT	: inout std_logic ;
			
		-- General Purpose I/O
		HPS_GPIO				: inout std_logic_vector(1 downto 0);
		
		-- I2C
		HPS_I2C_CONTROL	: inout std_logic ;
		HPS_I2C1_SCLK		: inout std_logic ;
		HPS_I2C1_SDAT		: inout std_logic ;
		HPS_I2C2_SCLK		: inout std_logic ;
		HPS_I2C2_SDAT		: inout std_logic ;
	
		-- Pushbutton
		HPS_KEY				: inout std_logic ;
	
		-- LED
		HPS_LED				: inout std_logic ;
			
		-- SD Card
		HPS_SD_CLK			: out std_logic ;
		HPS_SD_CMD			: inout std_logic ;
		HPS_SD_DATA			: inout std_logic_vector(3 downto 0) ;
	
		-- SPI
		HPS_SPIM_CLK		: out std_logic ;
		HPS_SPIM_MISO		: in std_logic ;
		HPS_SPIM_MOSI		: out std_logic ;
		HPS_SPIM_SS			: inout std_logic ;
	
		-- UART
		HPS_UART_RX			: in std_logic ;
		HPS_UART_TX			: out std_logic ;
	
		-- USB
		HPS_CONV_USB_N			: inout std_logic ;
		HPS_USB_CLKOUT			: in std_logic ;
		HPS_USB_DATA			: inout std_logic_vector(7 downto 0) ;
		HPS_USB_DIR				: in std_logic ;
		HPS_USB_NXT				: in std_logic ;
		HPS_USB_STP				: out std_logic  
	 ) ;
END ;		-- end of entity


Architecture RTL of MyComputer is
-------------------------------------------------------------------------------------------
--  signal declarations for temporary signals/wires to connect sub-systems together
-------------------------------------------------------------------------------------------

		-- temp signals carrying 2 sets of 4 bit data to each pair of Hex displays
		-- The 3 pairs of 8 bit ports generated by QSYS will drive these wires
		-- and they will be connected to the 7-Segment decoders created in VHDL 
		-- and they will drive the real HEX display on the DE1
		
		Signal	Temp_hex0_1 								: std_logic_vector(7 downto 0)	;
		Signal	Temp_hex2_3 								: std_logic_vector(7 downto 0)	;
		Signal	Temp_hex4_5 								: std_logic_vector(7 downto 0)	;
	 
	 
		-- TEMP SIGNALS TO CONNECT IO BRIDGE from QSYS generated IOBridge TO SUBSYSTEMS INCLUDING GRAPHICS AND IO DEVICE (RS232'S)
   
		SIGNAL 	IO_IRQ_WIRE                          :  std_logic;
		SIGNAL 	IO_Address_WIRE                      :  std_logic_vector(15 downto 0);                    
		SIGNAL 	IO_Bus_Enable_WIRE                   :  std_logic;                                        
		SIGNAL 	IO_Byte_Enable_WIRE                  :  std_logic_vector(1 downto 0);                     
		SIGNAL 	IO_RW_WIRE                           :  std_logic;                                        
		SIGNAL 	IO_Write_Data_WIRE                   :  std_logic_vector(15 downto 0);                    
		SIGNAL 	IO_Read_Data_WIRE                    :  std_logic_vector(15 downto 0);
		
		-- Other temporary signals 
		SIGNAL	RESET_L_WIRE 								 :  STD_LOGIC;
		SIGNAL	IO_Enable_L_WIRE 							 :  STD_LOGIC;
		SIGNAL	IO_UpperByte_Select_L_WIRE 			 :  STD_LOGIC;
		SIGNAL	IO_LowerByte_Select_L_WIRE 			 :  STD_LOGIC;
			 
	 ---------------------------------------------------------------------------------------
	 -- declaration of a System that we will build based on the QSys generated systems
	 ---------------------------------------------------------------------------------------

	component CPEN391_Computer is
        port (
				---------------------------------------------------------------------------------------------
				-- FPGA Side
				---------------------------------------------------------------------------------------------
				
				---------------------------------------------------------------------------------------------
				-- LEDS and Slider Switches
				---------------------------------------------------------------------------------------------
				leds_export                     : out   std_logic_vector(9 downto 0);
            slider_switches_export          : in    std_logic_vector(9 downto 0)  := (others => 'X');

				---------------------------------------------------------------------------------------------
				-- 7-Segment Displays
				-- These are the names of the exported 7-Segment display created in QSys
				---------------------------------------------------------------------------------------------
				hex0_1_export                   : out   std_logic_vector(7 downto 0);
				hex2_3_export                   : out   std_logic_vector(7 downto 0);
				hex4_5_export                   : out   std_logic_vector(7 downto 0);
				
				---------------------------------------------------------------------------------------------
				-- Push button
				---------------------------------------------------------------------------------------------
				pushbuttons_export              : in    std_logic_vector(3 downto 0)  := (others => 'X');
				
				-----------------------------------------------------------------------------
				-- LCD Exported Signals
				-----------------------------------------------------------------------------
				
				lcd_RS         						: out   std_logic;
				lcd_RW         						: out   std_logic;
				lcd_data       						: inout std_logic_vector(7 downto 0)  := (others => 'X');
				lcd_EN         						: out   std_logic;
				lcd_ON         						: out   std_logic;
				lcd_BLON       						: out   std_logic;
		
				-----------------------------------------------------------------------------
				-- Io Bridge Exported Signals
				-----------------------------------------------------------------------------
				io_acknowledge                  : in    std_logic                     := '0';             
				io_irq                          : in    std_logic                     := '0';             
				io_address                      : out   std_logic_vector(15 downto 0);                    
				io_bus_enable                   : out   std_logic;                                        
				io_byte_enable                  : out   std_logic_vector(1 downto 0);                     
				io_rw                           : out   std_logic;                                        
				io_write_data                   : out   std_logic_vector(15 downto 0);                    
				io_read_data                    : in    std_logic_vector(15 downto 0) := (others => '0');				
            
				---------------------------------------------------------------------------------------------
				-- SDRam on FPGA Side
				---------------------------------------------------------------------------------------------
				sdram_addr                      : out   std_logic_vector(12 downto 0);
            sdram_ba                        : out   std_logic_vector(1 downto 0);
            sdram_cas_n                     : out   std_logic;
            sdram_cke                       : out   std_logic;
            sdram_cs_n                      : out   std_logic;
            sdram_dq                        : inout std_logic_vector(15 downto 0) := (others => 'X');
            sdram_dqm                       : out   std_logic_vector(1 downto 0);
            sdram_ras_n                     : out   std_logic;
            sdram_we_n                      : out   std_logic;
            sdram_clk_clk                   : out   std_logic;
            
				---------------------------------------------------------------------------------------------
				-- HPS Side
				---------------------------------------------------------------------------------------------
				hps_io_hps_io_emac1_inst_TX_CLK : out   std_logic;
            hps_io_hps_io_emac1_inst_TXD0   : out   std_logic;
            hps_io_hps_io_emac1_inst_TXD1   : out   std_logic;
            hps_io_hps_io_emac1_inst_TXD2   : out   std_logic;
            hps_io_hps_io_emac1_inst_TXD3   : out   std_logic;
            hps_io_hps_io_emac1_inst_RXD0   : in    std_logic                     := 'X';
            hps_io_hps_io_emac1_inst_MDIO   : inout std_logic                     := 'X';
            hps_io_hps_io_emac1_inst_MDC    : out   std_logic;
            hps_io_hps_io_emac1_inst_RX_CTL : in    std_logic                     := 'X';
            hps_io_hps_io_emac1_inst_TX_CTL : out   std_logic;
            hps_io_hps_io_emac1_inst_RX_CLK : in    std_logic                     := 'X';
            hps_io_hps_io_emac1_inst_RXD1   : in    std_logic                     := 'X';
            hps_io_hps_io_emac1_inst_RXD2   : in    std_logic                     := 'X';
            hps_io_hps_io_emac1_inst_RXD3   : in    std_logic                     := 'X';
            hps_io_hps_io_qspi_inst_IO0     : inout std_logic                     := 'X';
            hps_io_hps_io_qspi_inst_IO1     : inout std_logic                     := 'X';
            hps_io_hps_io_qspi_inst_IO2     : inout std_logic                     := 'X';
            hps_io_hps_io_qspi_inst_IO3     : inout std_logic                     := 'X';
            hps_io_hps_io_qspi_inst_SS0     : out   std_logic;
            hps_io_hps_io_qspi_inst_CLK     : out   std_logic;
            hps_io_hps_io_sdio_inst_CMD     : inout std_logic                     := 'X';
            hps_io_hps_io_sdio_inst_D0      : inout std_logic                     := 'X';
            hps_io_hps_io_sdio_inst_D1      : inout std_logic                     := 'X';
            hps_io_hps_io_sdio_inst_CLK     : out   std_logic;
            hps_io_hps_io_sdio_inst_D2      : inout std_logic                     := 'X';
            hps_io_hps_io_sdio_inst_D3      : inout std_logic                     := 'X';
            hps_io_hps_io_usb1_inst_D0      : inout std_logic                     := 'X';
            hps_io_hps_io_usb1_inst_D1      : inout std_logic                     := 'X';
            hps_io_hps_io_usb1_inst_D2      : inout std_logic                     := 'X';
            hps_io_hps_io_usb1_inst_D3      : inout std_logic                     := 'X';
            hps_io_hps_io_usb1_inst_D4      : inout std_logic                     := 'X';
            hps_io_hps_io_usb1_inst_D5      : inout std_logic                     := 'X';
            hps_io_hps_io_usb1_inst_D6      : inout std_logic                     := 'X'; 
            hps_io_hps_io_usb1_inst_D7      : inout std_logic                     := 'X';
            hps_io_hps_io_usb1_inst_CLK     : in    std_logic                     := 'X';
            hps_io_hps_io_usb1_inst_STP     : out   std_logic;
            hps_io_hps_io_usb1_inst_DIR     : in    std_logic                     := 'X';
            hps_io_hps_io_usb1_inst_NXT     : in    std_logic                     := 'X';
            hps_io_hps_io_spim1_inst_CLK    : out   std_logic;
            hps_io_hps_io_spim1_inst_MOSI   : out   std_logic;
            hps_io_hps_io_spim1_inst_MISO   : in    std_logic                     := 'X';
            hps_io_hps_io_spim1_inst_SS0    : out   std_logic;
            hps_io_hps_io_uart0_inst_RX     : in    std_logic                     := 'X';
            hps_io_hps_io_uart0_inst_TX     : out   std_logic;
            hps_io_hps_io_i2c0_inst_SDA     : inout std_logic                     := 'X';
            hps_io_hps_io_i2c0_inst_SCL     : inout std_logic                     := 'X';
            hps_io_hps_io_i2c1_inst_SDA     : inout std_logic                     := 'X';
            hps_io_hps_io_i2c1_inst_SCL     : inout std_logic                     := 'X';
            hps_io_hps_io_gpio_inst_GPIO09  : inout std_logic                     := 'X';
            hps_io_hps_io_gpio_inst_GPIO35  : inout std_logic                     := 'X';
            hps_io_hps_io_gpio_inst_GPIO40  : inout std_logic                     := 'X';
            hps_io_hps_io_gpio_inst_GPIO41  : inout std_logic                     := 'X';
            hps_io_hps_io_gpio_inst_GPIO48  : inout std_logic                     := 'X';
            hps_io_hps_io_gpio_inst_GPIO53  : inout std_logic                     := 'X';
            hps_io_hps_io_gpio_inst_GPIO54  : inout std_logic                     := 'X';
            hps_io_hps_io_gpio_inst_GPIO61  : inout std_logic                     := 'X';
            
				memory_mem_a                    : out   std_logic_vector(14 downto 0);
            memory_mem_ba                   : out   std_logic_vector(2 downto 0);
            memory_mem_ck                   : out   std_logic;
            memory_mem_ck_n                 : out   std_logic;
            memory_mem_cke                  : out   std_logic;
            memory_mem_cs_n                 : out   std_logic;
            memory_mem_ras_n                : out   std_logic;
            memory_mem_cas_n                : out   std_logic;
            memory_mem_we_n                 : out   std_logic;
            memory_mem_reset_n              : out   std_logic;
            memory_mem_dq                   : inout std_logic_vector(31 downto 0) := (others => 'X');
            memory_mem_dqs                  : inout std_logic_vector(3 downto 0)  := (others => 'X');
            memory_mem_dqs_n                : inout std_logic_vector(3 downto 0)  := (others => 'X');
            memory_mem_odt                  : out   std_logic;
            memory_mem_dm                   : out   std_logic_vector(3 downto 0);
            memory_oct_rzqin                : in    std_logic                     := 'X';
            
            system_pll_ref_clk_clk          : in    std_logic                     := 'X';
            system_pll_ref_reset_reset      : in    std_logic                     := 'X'
       );
    end component CPEN391_Computer;
	 
	 ---------------------------------------------------------------------------------------
	 -- declaration of a component for a 4 bit to 7 segment decoder
	 ---------------------------------------------------------------------------------------
	 component HexTo7SegmentDisplay is
		Port (
				Input1 : in std_logic_vector(7 downto 0);
				
				Display1 : out std_logic_vector(6 downto 0) ;
				Display0 : out std_logic_vector(6 downto 0) 
		);
	 END component HexTo7SegmentDisplay;
	
	
	---------------------------------------------------------------------------------------
	 -- declaration of a component for a graphics controller
	---------------------------------------------------------------------------------------
	COMPONENT graphics_and_video_controller
		PORT( Reset_L : IN STD_LOGIC;
			 Clock_50Mhz : IN STD_LOGIC;
			 IOEnable_L : IN STD_LOGIC;
			 UpperByteSelect_L : IN STD_LOGIC;
			 LowerByteSelect_L : IN STD_LOGIC;
			 WriteEnable_L : IN STD_LOGIC;
			 GraphicsCS_L : IN STD_LOGIC;
			 Address : IN STD_LOGIC_VECTOR(15 DOWNTO 0);
			 DataIn : IN STD_LOGIC_VECTOR(15 DOWNTO 0);
		    DataOut : OUT STD_LOGIC_VECTOR(15 DOWNTO 0);
			 ----------------------------------------------
			 VGA_Clock : OUT STD_LOGIC;
			 VGA_HSync : OUT STD_LOGIC;
			 VGA_VSync : OUT STD_LOGIC;
			 VGA_Blanking : OUT STD_LOGIC;
			 VGA_Sync : OUT STD_LOGIC;
			 VGA_Blue : OUT STD_LOGIC_VECTOR(7 DOWNTO 0);
			 VGA_Green : OUT STD_LOGIC_VECTOR(7 DOWNTO 0);
			 VGA_Red : OUT STD_LOGIC_VECTOR(7 DOWNTO 0)
		);
	END COMPONENT;	
		
	 ---------------------------------------------------------------------------------------
	 -- declaration of a component for the serial ports
	 ---------------------------------------------------------------------------------------
	COMPONENT OnChipM68xxIO
		PORT(
			 Clock_50Mhz : IN STD_LOGIC;
			 IOSelect_H : IN STD_LOGIC;
			 ByteSelect_L : IN STD_LOGIC;
			 WE_L : IN STD_LOGIC;
			 Reset_L : IN STD_LOGIC;
			 Address : IN STD_LOGIC_VECTOR(15 DOWNTO 0);
			 DataIn : IN STD_LOGIC_VECTOR(7 DOWNTO 0);
			 ACIA_IRQ : OUT STD_LOGIC;
			 -------------------------------------------
			 RS232_RxData : IN STD_LOGIC ;
			 RS232_TxData : OUT STD_LOGIC ;
			 
			 GPS_RxData : IN STD_LOGIC;
			 GPS_TxData : OUT STD_LOGIC;
			 
			 BlueTooth_RxData : IN STD_LOGIC;
			 BlueTooth_TxData : OUT STD_LOGIC;
			 
			 TouchScreen_RxData : IN STD_LOGIC;
			 TouchScreen_TxData : OUT STD_LOGIC;
			 
			 DataOut : OUT STD_LOGIC_VECTOR(7 DOWNTO 0)
		);
	END COMPONENT;

	 
--------------------------------------------------------------------------------------------------
-- Start of the Architecture where we Instantiate components and connect them to real
-- Hardware on the DE1 or to temporary signals connecting building blocks/sub-system together
--------------------------------------------------------------------------------------------------
	 
BEGIN	 

		RESET_L_WIRE <= '1';	 
		GPIO_1(10) <= '0' ;								-- connect contrast pin on 24x2 LCD display to ground
		
		-- connections to wires on the top level
		IO_Enable_L_WIRE 						<= NOT(IO_bus_enable_WIRE);
		IO_UpperByte_Select_L_WIRE 		<= NOT(IO_byte_enable_WIRE(1));		
		IO_LowerByte_Select_L_WIRE 		<= NOT(IO_byte_enable_WIRE(0));		
		
	 ---------------------------------------------------------------------------------------
	 -- u0 is an instanace of the QSYS generated computer
	 -- map its IO ports as described below
	 ---------------------------------------------------------------------------------------
		
		u0 : component CPEN391_Computer
        port map (
 				leds_export                     => LEDR,                    --  Leds exported in QSYS wired directly to Red LEDS on DE1
				pushbuttons_export              => KEY,     						--  Pushbuttons exported in QSYS wired directly to push button switches on DE1, 
																								--  thus, combined with settings when we created with QSYS makes give them interrupts capability
																								--  when pressed
				slider_switches_export          => SW,          				--  Slider_switches exported in QSYS wired directly to Slider switches on DE1

				-- port map, wire the exported QSYS generated 8 bit ports to temporary wires/signals
				hex0_1_export    							=> Temp_hex0_1,
            hex2_3_export    							=> Temp_hex2_3,
            hex4_5_export    							=> Temp_hex4_5,
				
				-- port map for the IO Bridge to temporary wires
				io_acknowledge  							=> IO_Bus_Enable_WIRE,	-- connect enable back to into acknowledge
				io_irq          							=> IO_IRQ_WIRE,
				io_address      							=> IO_Address_WIRE,
				io_bus_enable  							=> IO_Bus_Enable_WIRE,
				io_byte_enable  							=> IO_Byte_Enable_WIRE,
				io_rw           							=> IO_RW_WIRE,  
				io_write_data   							=> IO_Write_Data_WIRE,                    
				io_read_data    							=> IO_Read_Data_WIRE,
				
				-- Connect QSYS generated LCD display to the GPIO Pins
				lcd_DATA(0)    							=> GPIO_1(0),
				lcd_DATA(1)    							=> GPIO_1(1),
				lcd_DATA(2)    							=> GPIO_1(2),
				lcd_DATA(3)    							=> GPIO_1(3),
				lcd_DATA(4)   								=> GPIO_1(4),
				lcd_DATA(5)    							=> GPIO_1(5),
				lcd_DATA(6)    							=> GPIO_1(6),
				lcd_DATA(7)    							=> GPIO_1(7),

				-- lcd_ON         -- no connection on the actual 24 x 2 LCD display
				-- lcd_BLON       -- no connection on the actual 24 x 2 LCD display
				
				lcd_EN         							=> GPIO_1(13),
				lcd_RS        								=> GPIO_1(11),
				lcd_RW         							=> GPIO_1(15),
  
				-- port map, wire the exported QSYS generated SDRAM port directly to SDRAM chips on FPGA
				sdram_addr                      		=> DRAM_ADDR, 
            sdram_ba                       		=> DRAM_BA,
            sdram_cas_n                    	 	=> DRAM_CAS_N,
            sdram_cke                       		=> DRAM_CKE,
            sdram_cs_n                      		=> DRAM_CS_N,
            sdram_dq                        		=> DRAM_DQ,
            sdram_dqm(1)                    		=> DRAM_UDQM, 
				sdram_dqm(0)						  		=> DRAM_LDQM, 
            sdram_ras_n                     		=> DRAM_RAS_N,
            sdram_we_n                     		=> DRAM_WE_N,
            sdram_clk_clk	                 		=> DRAM_CLK,
           
 				-- port map, wire the exported ARM Cores (HPS) signals to PINs on DE1               
				hps_io_hps_io_emac1_inst_TX_CLK => HPS_ENET_GTX_CLK, 	
            hps_io_hps_io_emac1_inst_TXD0   => HPS_ENET_TX_DATA(0), 
            hps_io_hps_io_emac1_inst_TXD1   => HPS_ENET_TX_DATA(1),
            hps_io_hps_io_emac1_inst_TXD2   => HPS_ENET_TX_DATA(2),
            hps_io_hps_io_emac1_inst_TXD3   => HPS_ENET_TX_DATA(3),
            hps_io_hps_io_emac1_inst_RXD0   => HPS_ENET_RX_DATA(0), 
            hps_io_hps_io_emac1_inst_MDIO   => HPS_ENET_MDIO, 
            hps_io_hps_io_emac1_inst_MDC    => HPS_ENET_MDC,
            hps_io_hps_io_emac1_inst_RX_CTL => HPS_ENET_RX_DV, 
            hps_io_hps_io_emac1_inst_TX_CTL => HPS_ENET_TX_EN, 
            hps_io_hps_io_emac1_inst_RX_CLK => HPS_ENET_RX_CLK, 
            hps_io_hps_io_emac1_inst_RXD1   => HPS_ENET_RX_DATA(1),
            hps_io_hps_io_emac1_inst_RXD2   => HPS_ENET_RX_DATA(2), 
            hps_io_hps_io_emac1_inst_RXD3   => HPS_ENET_RX_DATA(3),
            hps_io_hps_io_qspi_inst_IO0     => HPS_FLASH_DATA(0), 
            hps_io_hps_io_qspi_inst_IO1     => HPS_FLASH_DATA(1),
            hps_io_hps_io_qspi_inst_IO2     => HPS_FLASH_DATA(2),
            hps_io_hps_io_qspi_inst_IO3     => HPS_FLASH_DATA(3),
            hps_io_hps_io_qspi_inst_SS0     => HPS_FLASH_NCSO,  
            hps_io_hps_io_qspi_inst_CLK     => HPS_FLASH_DCLK,
            hps_io_hps_io_sdio_inst_CMD     => HPS_SD_CMD,
            hps_io_hps_io_sdio_inst_D0      => HPS_SD_DATA(0),
            hps_io_hps_io_sdio_inst_D1      => HPS_SD_DATA(1),
            hps_io_hps_io_sdio_inst_CLK     => HPS_SD_CLK,
            hps_io_hps_io_sdio_inst_D2      => HPS_SD_DATA(2),
            hps_io_hps_io_sdio_inst_D3      => HPS_SD_DATA(3),
            hps_io_hps_io_usb1_inst_D0      => HPS_USB_DATA(0),
            hps_io_hps_io_usb1_inst_D1      => HPS_USB_DATA(1),
            hps_io_hps_io_usb1_inst_D2      => HPS_USB_DATA(2),
            hps_io_hps_io_usb1_inst_D3      => HPS_USB_DATA(3),
            hps_io_hps_io_usb1_inst_D4      => HPS_USB_DATA(4),
            hps_io_hps_io_usb1_inst_D5      => HPS_USB_DATA(5),
            hps_io_hps_io_usb1_inst_D6      => HPS_USB_DATA(6),
            hps_io_hps_io_usb1_inst_D7      => HPS_USB_DATA(7),
            hps_io_hps_io_usb1_inst_CLK     => HPS_USB_CLKOUT,
            hps_io_hps_io_usb1_inst_STP     => HPS_USB_STP,
            hps_io_hps_io_usb1_inst_DIR     => HPS_USB_DIR, 
            hps_io_hps_io_usb1_inst_NXT     => HPS_USB_NXT,
            hps_io_hps_io_spim1_inst_CLK    => HPS_SPIM_CLK,
            hps_io_hps_io_spim1_inst_MOSI   => HPS_SPIM_MOSI,
            hps_io_hps_io_spim1_inst_MISO   => HPS_SPIM_MISO,
            hps_io_hps_io_spim1_inst_SS0    => HPS_SPIM_SS, 
            hps_io_hps_io_uart0_inst_RX     => HPS_UART_RX,
            hps_io_hps_io_uart0_inst_TX     => HPS_UART_TX,
            hps_io_hps_io_i2c0_inst_SDA     => HPS_I2C1_SDAT,
            hps_io_hps_io_i2c0_inst_SCL     => HPS_I2C1_SCLK,
            hps_io_hps_io_i2c1_inst_SDA     => HPS_I2C2_SDAT, 
            hps_io_hps_io_i2c1_inst_SCL     => HPS_I2C2_SCLK,
            hps_io_hps_io_gpio_inst_GPIO09  => HPS_CONV_USB_N, 
            hps_io_hps_io_gpio_inst_GPIO35  => HPS_ENET_INT_N, 
            hps_io_hps_io_gpio_inst_GPIO40  => HPS_GPIO(0), 
            hps_io_hps_io_gpio_inst_GPIO41  => HPS_GPIO(1), 
            hps_io_hps_io_gpio_inst_GPIO48  => HPS_I2C_CONTROL, 
            hps_io_hps_io_gpio_inst_GPIO53  => HPS_LED,
            hps_io_hps_io_gpio_inst_GPIO54  => HPS_KEY,
            hps_io_hps_io_gpio_inst_GPIO61  => HPS_GSENSOR_INT,
            
				memory_mem_a                    => HPS_DDR3_ADDR,
            memory_mem_ba                   => HPS_DDR3_BA,
            memory_mem_ck                   => HPS_DDR3_CK_P,
            memory_mem_ck_n                 => HPS_DDR3_CK_N,
            memory_mem_cke                  => HPS_DDR3_CKE, 
            memory_mem_cs_n                 => HPS_DDR3_CS_N,
            memory_mem_ras_n                => HPS_DDR3_RAS_N,
            memory_mem_cas_n                => HPS_DDR3_CAS_N,
            memory_mem_we_n                 => HPS_DDR3_WE_N,
            memory_mem_reset_n              => HPS_DDR3_RESET_N,
            memory_mem_dq                   => HPS_DDR3_DQ,
            memory_mem_dqs                  => HPS_DDR3_DQS_P,
            memory_mem_dqs_n                => HPS_DDR3_DQS_N,
            memory_mem_odt                  => HPS_DDR3_ODT,
            memory_mem_dm                   => HPS_DDR3_DM,
            memory_oct_rzqin                => HPS_DDR3_RZQ,
				
				system_pll_ref_clk_clk          => CLOCK_50, 
            system_pll_ref_reset_reset      => '0'
        );
		  
		  -----------------------------------------------------------------------------------------------
		  -- Instantiate 3 instances of the seven seg decoders
		  -- one for hex display 0 and 1
		  -- one for hex display 2 and 3
		  -- one for hex display 4 and 5
		  -- Connect their inputs to the temporary wires/signals being driven by the ports
		  -- exported in Qsys and connect their outputs to the real 7-Segment displays on the DE1
		  -----------------------------------------------------------------------------------------------
		  
		  HEXDisplay0_1 : component HexTo7SegmentDisplay			-- HEXDisplay0_1 is an instance of pair of 7 segment decoder
				Port Map (
						-- inputs
						Input1 => Temp_hex0_1,								-- Connect input1 of the HexDisplay circuit to temporary signal/wire

						-- outputs: Mapping important
						Display0(6 downto 0) => HEX0(6 downto 0),		-- output of the component connect to HEX displays 0 and 1 on the DE1
						Display1(6 downto 0) => HEX1(6 downto 0)		-- output of the component connect to HEX displays 0 and 1 on the DE1
				);
				
			HEXDisplay2_3 : component HexTo7SegmentDisplay			-- HEXDisplay2_3 is an instance of pair of 7 segment decoder
				Port Map (
						-- inputs
						Input1 => Temp_hex2_3,								-- Connect input1 of the HexDisplay circuit to temporary signal/wire

						-- outputs: Mapping important
						Display0(6 downto 0) => HEX2(6 downto 0),		-- output of the component connect to HEX displays 2 and 3 on the DE1
						Display1(6 downto 0) => HEX3(6 downto 0)		-- output of the component connect to HEX displays 2 and 3 on the DE1
				);
				
		  HEXDisplay4_5 : component HexTo7SegmentDisplay			-- HEXDisplay4_5 is an instance of pair of 7 segment decoder
				Port Map (
						-- inputs
						Input1 => Temp_hex4_5,								-- Connect input1 of the HexDisplay circuit to temporary signal/wire

						-- outputs: Mapping important
						Display0(6 downto 0) => HEX4(6 downto 0),		-- output of the component connect to HEX displays 4 and 5 on the DE1
						Display1(6 downto 0) => HEX5(6 downto 0)		-- output of the component connect to HEX displays 4 and 5 on the DE1
				);
			
		-- create an instance of the graphics controller
		GraphicsController1 : graphics_and_video_controller
			PORT MAP(
				Reset_L 							=> Reset_L_WIRE,
				Clock_50Mhz 					=> CLOCK_50,
				Address 							=> IO_Address_WIRE,
				DataIn 							=> IO_Write_Data_WIRE,
				DataOut 							=> IO_Read_Data_WIRE,
				IOEnable_L 						=> IO_Enable_L_WIRE,
				UpperByteSelect_L 			=> IO_UpperByte_Select_L_WIRE,
				LowerByteSelect_L 			=> IO_LowerByte_Select_L_WIRE,
				WriteEnable_L 					=> IO_RW_WIRE,
				GraphicsCS_L 					=> IO_Enable_L_WIRE,
				--
				VGA_Clock						=> VGA_Clk,
				VGA_Blue 						=> VGA_B,
				VGA_Green 						=> VGA_G,
				VGA_Red							=> VGA_R,
				VGA_HSync 						=> VGA_HS,
				VGA_VSync						=> VGA_VS,
				VGA_Blanking 					=> VGA_BLANK_N,
				VGA_SYNC							=> VGA_SYNC_N
		 );	
		 
		-- create an instance of the IO port with serial ports
		
		 IOPorts : OnChipM68xxIO
			 PORT MAP(
				 -- Bridge Signals
				 Reset_L 									=> Reset_L_WIRE,
				 Clock_50Mhz 								=> CLOCK_50,
				 Address 									=> IO_Address_WIRE,
				 DataIn 										=> IO_Write_Data_WIRE(7 DOWNTO 0),
				 DataOut 									=> IO_Read_Data_WIRE(7 DOWNTO 0),
				 IOSelect_H 								=> IO_Bus_Enable_WIRE,
				 ByteSelect_L 								=> IO_LowerByte_Select_L_WIRE,
				 WE_L 										=> IO_RW_WIRE,
				 ACIA_IRQ 									=> IO_IRQ_WIRE,
				 
				 -- Real World Signals
				 RS232_RxData								=> GPIO_1(29),
				 RS232_TxData								=> GPIO_1(27),

				 GPS_RxData 								=> GPIO_1(28),
				 GPS_TxData 								=> GPIO_1(26),

				 BlueTooth_RxData 						=> GPIO_1(18),
				 BlueTooth_TxData 						=> GPIO_1(19),
				 
				 TouchScreen_RxData 						=> GPIO_0(11),
				 TouchScreen_TxData 						=> GPIO_0(10)
		);
end ;
